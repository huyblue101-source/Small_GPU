module top (
    input wire clk,
    input wire reset
);

// TODO: connect GPU modules here

endmodule
